library verilog;
use verilog.vl_types.all;
entity ALU1BIT_vlg_vec_tst is
end ALU1BIT_vlg_vec_tst;
