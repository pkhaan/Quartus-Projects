library verilog;
use verilog.vl_types.all;
entity Problem1_vlg_vec_tst is
end Problem1_vlg_vec_tst;
