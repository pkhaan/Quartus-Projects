library verilog;
use verilog.vl_types.all;
entity ERG1PR3_vlg_check_tst is
    port(
        f               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end ERG1PR3_vlg_check_tst;
