library verilog;
use verilog.vl_types.all;
entity ALU16BIT_vlg_vec_tst is
end ALU16BIT_vlg_vec_tst;
