library verilog;
use verilog.vl_types.all;
entity Lab1b_vlg_vec_tst is
end Lab1b_vlg_vec_tst;
