library verilog;
use verilog.vl_types.all;
entity Problem1_vlg_check_tst is
    port(
        f               : in     vl_logic;
        g               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end Problem1_vlg_check_tst;
