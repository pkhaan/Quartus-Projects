library verilog;
use verilog.vl_types.all;
entity ask2_vlg_check_tst is
    port(
        f               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end ask2_vlg_check_tst;
