LIBRARY ieee ;
USE ieee.std_logic_1164.all ;
USE ieee.std_logic_signed.all ;

ENTITY vend IS
	PORT ( N, D, Q, Resetn, Coin : IN STD_LOGIC ;
		 Z 			     : OUT STD_LOGIC ) ;
END vend ;

ARCHITECTURE Behavior OF vend IS
	SIGNAL X: STD_LOGIC_VECTOR(4 DOWNTO 0) ;
	SIGNAL S: STD_LOGIC_VECTOR(5 DOWNTO 0) ;
BEGIN
	X(0) <= N OR Q ;
	X(1) <= D ;
	X(2) <= N ;
	X(3) <= D OR Q ;
	X(4) <= Q ;
	PROCESS ( Resetn, Coin )
	BEGIN
		IF Resetn = '0' THEN
			S <= "000000" ;
		ELSIF Coin'EVENT AND Coin = '0' THEN
			S <= ('0' & X) + S ;
		END IF ;
	END PROCESS ;
	Z <= S(5) OR (S(4) AND S(3) AND S(2) AND S(1)) ;
END Behavior ;