library verilog;
use verilog.vl_types.all;
entity ERG1PR3_vlg_vec_tst is
end ERG1PR3_vlg_vec_tst;
