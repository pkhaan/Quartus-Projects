library verilog;
use verilog.vl_types.all;
entity Problem2_vlg_vec_tst is
end Problem2_vlg_vec_tst;
