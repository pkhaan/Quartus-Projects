library verilog;
use verilog.vl_types.all;
entity Problem2 is
    port(
        f               : out    vl_logic;
        x2              : in     vl_logic;
        x1              : in     vl_logic;
        x4              : in     vl_logic;
        x3              : in     vl_logic
    );
end Problem2;
