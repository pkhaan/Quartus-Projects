library verilog;
use verilog.vl_types.all;
entity ask2_vlg_vec_tst is
end ask2_vlg_vec_tst;
