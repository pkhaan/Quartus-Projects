library verilog;
use verilog.vl_types.all;
entity VHDLEXAMPLE_vlg_vec_tst is
end VHDLEXAMPLE_vlg_vec_tst;
