library verilog;
use verilog.vl_types.all;
entity ERGASTHRIO1_vlg_vec_tst is
end ERGASTHRIO1_vlg_vec_tst;
