library verilog;
use verilog.vl_types.all;
entity Problem1 is
    port(
        x1              : in     vl_logic;
        x2              : in     vl_logic;
        x3              : in     vl_logic;
        x4              : in     vl_logic;
        x5              : in     vl_logic;
        f               : out    vl_logic;
        g               : out    vl_logic
    );
end Problem1;
